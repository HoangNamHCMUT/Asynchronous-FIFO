
`define PTR_WIDTH 4

`define WIDTH 4
